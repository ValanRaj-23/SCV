module()
endmodule
